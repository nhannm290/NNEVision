module Convolution_layer1 (
    input [31:0] Data_In
);
    
endmodule