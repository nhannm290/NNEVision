module Sigmol (
    input [31:0] Data_In,
    input clk,
    input rst,
    input Valid_In,
    output [31:0] Data_Out,
    output Valid_Out
);
    
endmodule