module Kernel_3x3_stride_1x1 (
    ports
);
    
endmodule