module Test_Convolution2D_3x3_stride_1x1_padding_1x1 (
    
);
    parameter DATA_WIDHT = 32;
    parameter IMG_WIDHT = 220;
    parameter   IMG_HEIGHT =220;

    
    
endmodule