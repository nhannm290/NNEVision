module Layer2 #(
    parameter DATA_WIDHT = 32,
    parameter IMG_WIDHT =220,
    parameter IMG_HEIGHT =220
) (
    input [DATA_WIDHT*8-1:0] Data_In,
    input clk,
    input rst,
    input Valid_In,
    output [DATA_WIDHT*8-1:0] Data_Out1,
    output Valid_Out 
);


    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL1_K1(
            .Data_In(Data_In[DATA_WIDHT-1:0]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );

    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL2_K1(
            .Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );

    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL3_K1(
            .Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );

    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL4_K1(
            .Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );

    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL5_K1(
            .Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );

    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL6_K1(
            .Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );
    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL7_K1(
            .Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );    

    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL8_K1(
            .Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );
    ///////////////////////// KERNEL 2
    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL1_K(
            .Data_In(Data_In[DATA_WIDHT-1:0]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );

    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL2_1(
            .Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );

    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL3_K1(
            .Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );

    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL4_K1(
            .Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );

    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL5_K1(
            .Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );

    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL6_K1(
            .Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );
    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL7_K1(
            .Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );    

    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL8_K1(
            .Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );
/////////////////////////////// KERNEL 3
    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL1_K1(
            .Data_In(Data_In[DATA_WIDHT-1:0]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );

    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL2_1(
            .Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );

    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL3_K1(
            .Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );

    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL4_K1(
            .Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );

    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL5_K1(
            .Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );

    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL6_K1(
            .Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );
    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL7_K1(
            .Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );    

    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL8_K1(
            .Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );
////////////////////////////// KERNEL 4
    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL1_K1(
            .Data_In(Data_In[DATA_WIDHT-1:0]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );

    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL2_1(
            .Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );

    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL3_K1(
            .Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );

    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL4_K1(
            .Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );

    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL5_K1(
            .Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );

    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL6_K1(
            .Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );
    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL7_K1(
            .Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );    

    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL8_K1(
            .Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );
//////////////////////// Kernel 5
    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL1_K1(
            .Data_In(Data_In[DATA_WIDHT-1:0]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );

    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL2_1(
            .Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );

    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL3_K1(
            .Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );

    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL4_K1(
            .Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );

    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL5_K1(
            .Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );

    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL6_K1(
            .Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );
    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL7_K1(
            .Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );    

    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL8_K1(
            .Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );
//////////////////////////////////// KERNEl 6
    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL1_K1(
            .Data_In(Data_In[DATA_WIDHT-1:0]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );

    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL2_1(
            .Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );

    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL3_K1(
            .Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );

    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL4_K1(
            .Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );

    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL5_K1(
            .Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );

    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL6_K1(
            .Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );
    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL7_K1(
            .Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );    

    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL8_K1(
            .Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );
//////////////////////////////// KERNEL 7
    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL1_K1(
            .Data_In(Data_In[DATA_WIDHT-1:0]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );

    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL2_1(
            .Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );

    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL3_K1(
            .Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );

    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL4_K1(
            .Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );

    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL5_K1(
            .Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );

    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL6_K1(
            .Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );
    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL7_K1(
            .Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );    

    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL8_K1(
            .Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );
////////////////////////////////// KERNEL 8
    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL1_K1(
            .Data_In(Data_In[DATA_WIDHT-1:0]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );

    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL2_1(
            .Data_In(Data_In[DATA_WIDHT*2-1:DATA_WIDHT]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );

    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL3_K1(
            .Data_In(Data_In[DATA_WIDHT*3-1:DATA_WIDHT*2]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );

    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL4_K1(
            .Data_In(Data_In[DATA_WIDHT*4-1:DATA_WIDHT*3]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );

    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL5_K1(
            .Data_In(Data_In[DATA_WIDHT*5-1:DATA_WIDHT*4]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );

    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL6_K1(
            .Data_In(Data_In[DATA_WIDHT*6-1:DATA_WIDHT*5]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );
    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL7_K1(
            .Data_In(Data_In[DATA_WIDHT*7-1:DATA_WIDHT*6]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );    

    Covolution2D_3x3_stride1x1 #(
        .DATA_WIDHT(DATA_WIDHT),
        .IMG_WIDTH(IMG_WIDTH),
        .IMG_HEIGHT(IMG_HEIGHT),
        )
        CHANNEL8_K1(
            .Data_In(Data_In[DATA_WIDHT*8-1:DATA_WIDHT*7]),
            .Kernel1({}),
            .Kernel2(0),
            .Kernel3(0),
            .Kernel4(0),
            .Kernel5(0),
            .Kernel6(0),
            .Kernel7(0),
            .Kernel8(0),
            .Kernel9(0),
            .clk(clk),
            .rst(rst),
            .Valid_In(Valid_In),
            .Data_Out(),
            .Valid_Out()
        );                

endmodule